package test_pkg;
	
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "src_agent_config.sv"
	`include "dst_agent_config.sv"
	`include "env_config.sv"
	`include "src_xtn.sv"

	`include "src_driver.sv"
	`include "src_monitor.sv"
	`include "src_sequencer.sv"
	`include "src_agent.sv"
	`include "src_agent_top.sv"
	//`include "src_seqs.sv"

	`include "dst_xtn.sv"
	`include "dst_monitor.sv"
	`include "dst_sequencer.sv"
	//`include "dst_seqs.sv"
	`include "dst_driver.sv"
	`include "dst_agent.sv"
	`include "dst_agent_top.sv"

	//`include "ram_virtual_sequencer.sv"
	//`include "ram_virtual_seqs.sv"
	`include "scoreboard.sv"

	`include "tb.sv"


	`include "vtest_lib.sv"
	
endpackage
