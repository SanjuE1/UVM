class src_xtn extends uvm_sequence_item;
	`uvm_object_utils(src_xtn)
	function new(string name="src_xtn");
		super.new(name);
	endfunction
endclass


