module top;
	
	import test_pkg::*;	
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	initial begin 
		run_test();
		end
endmodule

